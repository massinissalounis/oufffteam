-- Oufffteam
-- Projet carte m�re
-- Device: Debug PMP

-- 25/01/2010			CBE			Cr�ation

entity debug_pmp is

end entity debug_pmp;