-- Auteur: P.P
-- Version: A
-- Date de cr�ation: 12/01/11

-- Description: Top level entity du CPLD de la balise Rx
-- Cible: XC2C128 - VQ100

LIBRARY IEEE;
	USE IEEE.STD_LOGIC_1164.ALL;
	USE IEEE.NUMERIC_STD.ALL;

ENTITY RX_cpld IS
	PORT		(	-- I/O G�n�riques
					CLK		: IN STD_LOGIC;
					LED1		: OUT STD_LOGIC;
					LED2		: OUT STD_LOGIC;
					-- TSOPs
					TSOP1		: IN STD_LOGIC_VECTOR (15 DOWNTO 0);
					TSOP2		: IN STD_LOGIC_VECTOR (15 DOWNTO 0);
					-- PIC
					PIC_Rx		: OUT STD_LOGIC; -- PIC_CPLD PORT 9 USED AS SERIAL LINE (PIC's PIN36 - RP19)
					ADR			: IN STD_LOGIC_VECTOR (8 DOWNTO 0)); -- selection d'adresses pour les TSOP
END ENTITY RX_cpld;


ARCHITECTURE basic_mux_RX_cpld OF RX_cpld IS
SIGNAL INT_TSOP : STD_LOGIC_VECTOR (31 DOWNTO 0);
SIGNAL INT_ADR : STD_LOGIC_VECTOR (8 DOWNTO 0);
SIGNAL INT_PIC_Rx : STD_LOGIC;

BEGIN
	
	-- Assignation des signaux
	INT_TSOP(31 DOWNTO 16) <= TSOP1;
	INT_TSOP(15 DOWNTO 0) <= TSOP2;
	INT_ADR<=ADR;
	PIC_Rx <= INT_PIC_Rx;
	LED1 <= '1';
	LED2 <= NOT INT_PIC_Rx;
	
	--MUX
	WITH INT_ADR SELECT
		INT_PIC_Rx <=	INT_TSOP(0) WHEN "000000000",
							INT_TSOP(1) WHEN "000000001",
							INT_TSOP(2) WHEN "000000010",
							INT_TSOP(3) WHEN "000000011",
							INT_TSOP(4) WHEN "000000100",
							INT_TSOP(5) WHEN "000000101",
							INT_TSOP(6) WHEN "000000110",
							INT_TSOP(7) WHEN "000000111",
							INT_TSOP(8) WHEN "000001000",
							INT_TSOP(9) WHEN "000001001",
							INT_TSOP(10) WHEN "000001010",
							INT_TSOP(11) WHEN "000001011",
							INT_TSOP(12) WHEN "000001100",
							INT_TSOP(13) WHEN "000001101",
							INT_TSOP(14) WHEN "000001110",
							INT_TSOP(15) WHEN "000001111",
							INT_TSOP(16) WHEN "000010000",
							INT_TSOP(17) WHEN "000010001",
							INT_TSOP(18) WHEN "000010010",
							INT_TSOP(19) WHEN "000010011",
							INT_TSOP(20) WHEN "000010100",
							INT_TSOP(21) WHEN "000010101",
							INT_TSOP(22) WHEN "000010110",
							INT_TSOP(23) WHEN "000010111",
							INT_TSOP(24) WHEN "000011000",
							INT_TSOP(25) WHEN "000011001",
							INT_TSOP(26) WHEN "000011010",
							INT_TSOP(27) WHEN "000011011",
							INT_TSOP(28) WHEN "000011100",
							INT_TSOP(29) WHEN "000011101",
							INT_TSOP(30) WHEN "000011110",
							INT_TSOP(31) WHEN "000011111",
							'1' WHEN OTHERS;
END ARCHITECTURE;